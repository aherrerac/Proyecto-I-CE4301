module alu32(input logic [31:0] A, B,
 				 input logic [2:0] F,
				 output logic [31:0] Y,
				 output logic Negative, Zero, Carry,Overflow);
	logic [31:0] S, Bout;
	logic Cout;
	assign Bout = F[2] ? ~B : B;
	
	
	//assign S = A + Bout + F[2];
	
	//full_adder sum (A,Bout,F[2], S, Cout);
	assign {Cout, S} = A +Bout + F[2];
	
	
	always_comb
		case (F[1:0])
			2'b00: Y <= A & Bout;
			2'b01: Y <= A | Bout;
			2'b10: Y <= S;
			2'b11: Y <= S[31];
		endcase

	assign Zero = (Y == 0);
	assign Negative = (Y[31]==32'b1);
	/*assign Overflow = ~F[2] & (A & B & ~S[31] | ~A & ~B & S[31]) |
							 F[2] & (~A & B & S[31] | A & ~B & ~S[31]);*/
	always_comb
		case (F[2:1])
			2'b01: Overflow <= A[31] & (B[31] & ~S[31] | ~A[31] & ~B[31] & S[31]);
			2'b11: Overflow <= ~A[31] & (B[31] & S[31] | A[31] & ~B[31] & ~S[31]);
		default: Overflow <= 1'b0;
	endcase

	always_comb
		case (F[1:0])
			2'b10: Carry <= Cout;
			2'b11: Carry <= Cout;
		default: Carry <= 1'b0;
	endcase
	
endmodule