    Mac OS X            	   2   �      �                                      ATTR       �   �   %                  �   %  com.apple.quarantine q/0082;5be878a2;Telegram\x20Desktop; 