    Mac OS X            	   2   �      �                                      ATTR       �   �   5                  �     com.apple.lastuseddate#PS       �   %  com.apple.quarantine <��[    �}q    q/0082;5be8789e;Telegram\x20Desktop; 