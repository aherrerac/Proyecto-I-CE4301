    Mac OS X            	   2   �      �                                      ATTR       �   �   %                  �   %  com.apple.quarantine q/0082;5be878a1;Telegram\x20Desktop; 